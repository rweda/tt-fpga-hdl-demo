

// =======================
// The Tiny Tapeout module
// =======================

module tt_um_template (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    /*   // The FPGA is based on TinyTapeout 3 which has no bidirectional I/Os (vs. TT6 for the ASIC).
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    */
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
   logic passed, failed;  // Connected to uo_out[0] and uo_out[1] respectively, which connect to Makerchip passed/failed.

   wire reset = ! rst_n;

// ---------- Generated Code Inlined Here (before 1st \TLV) ----------
// Generated by SandPiper(TM) 1.14-2022/10/10-beta-Pro from Redwood EDA, LLC.
// (Installed here: /usr/local/mono/sandpiper/distro.)
// Redwood EDA, LLC does not claim intellectual property rights to this file and provides no warranty regarding its correctness or quality.


// For silencing unused signal messages.
`define BOGUS_USE(ignore)


genvar digit, dmem, imem, input_label, leds, switch, xreg;


//
// Signals declared top-level.
//

// For $slideswitch.
logic [7:0] L0_slideswitch_a0;

// For $sseg_decimal_point_n.
logic L0_sseg_decimal_point_n_a0;

// For $sseg_digit_n.
logic [7:0] L0_sseg_digit_n_a0;

// For $sseg_segment_n.
logic [6:0] L0_sseg_segment_n_a0;

// For /fpga_pins/fpga|cpu$br_tgt_pc.
logic [31:0] FpgaPins_Fpga_CPU_br_tgt_pc_a2,
             FpgaPins_Fpga_CPU_br_tgt_pc_a3;

// For /fpga_pins/fpga|cpu$dec_bits.
logic [10:0] FpgaPins_Fpga_CPU_dec_bits_a1;

// For /fpga_pins/fpga|cpu$dmem_addr.
logic [2:0] FpgaPins_Fpga_CPU_dmem_addr_a4;

// For /fpga_pins/fpga|cpu$dmem_rd_data.
logic [31:0] FpgaPins_Fpga_CPU_dmem_rd_data_a4,
             FpgaPins_Fpga_CPU_dmem_rd_data_a5;

// For /fpga_pins/fpga|cpu$dmem_rd_en.
logic FpgaPins_Fpga_CPU_dmem_rd_en_a4;

// For /fpga_pins/fpga|cpu$dmem_wr_data.
logic [31:0] FpgaPins_Fpga_CPU_dmem_wr_data_a4;

// For /fpga_pins/fpga|cpu$dmem_wr_en.
logic FpgaPins_Fpga_CPU_dmem_wr_en_a4;

// For /fpga_pins/fpga|cpu$funct3.
logic [2:0] FpgaPins_Fpga_CPU_funct3_a1;

// For /fpga_pins/fpga|cpu$funct3_valid.
logic FpgaPins_Fpga_CPU_funct3_valid_a1;

// For /fpga_pins/fpga|cpu$funct7.
logic [6:0] FpgaPins_Fpga_CPU_funct7_a1;

// For /fpga_pins/fpga|cpu$funct7_valid.
logic FpgaPins_Fpga_CPU_funct7_valid_a1;

// For /fpga_pins/fpga|cpu$imem_rd_addr.
logic [4-1:0] FpgaPins_Fpga_CPU_imem_rd_addr_a0,
              FpgaPins_Fpga_CPU_imem_rd_addr_a1;

// For /fpga_pins/fpga|cpu$imem_rd_data.
logic [31:0] FpgaPins_Fpga_CPU_imem_rd_data_a1;

// For /fpga_pins/fpga|cpu$imem_rd_en.
logic FpgaPins_Fpga_CPU_imem_rd_en_a0,
      FpgaPins_Fpga_CPU_imem_rd_en_a1;

// For /fpga_pins/fpga|cpu$imm.
logic [31:0] FpgaPins_Fpga_CPU_imm_a1,
             FpgaPins_Fpga_CPU_imm_a2,
             FpgaPins_Fpga_CPU_imm_a3;

// For /fpga_pins/fpga|cpu$inc_pc.
logic [31:0] FpgaPins_Fpga_CPU_inc_pc_a1,
             FpgaPins_Fpga_CPU_inc_pc_a2,
             FpgaPins_Fpga_CPU_inc_pc_a3;

// For /fpga_pins/fpga|cpu$instr.
logic [31:0] FpgaPins_Fpga_CPU_instr_a1;

// For /fpga_pins/fpga|cpu$is_add.
logic FpgaPins_Fpga_CPU_is_add_a1,
      FpgaPins_Fpga_CPU_is_add_a2,
      FpgaPins_Fpga_CPU_is_add_a3;

// For /fpga_pins/fpga|cpu$is_addi.
logic FpgaPins_Fpga_CPU_is_addi_a1,
      FpgaPins_Fpga_CPU_is_addi_a2,
      FpgaPins_Fpga_CPU_is_addi_a3;

// For /fpga_pins/fpga|cpu$is_and.
logic FpgaPins_Fpga_CPU_is_and_a1,
      FpgaPins_Fpga_CPU_is_and_a2,
      FpgaPins_Fpga_CPU_is_and_a3;

// For /fpga_pins/fpga|cpu$is_andi.
logic FpgaPins_Fpga_CPU_is_andi_a1,
      FpgaPins_Fpga_CPU_is_andi_a2,
      FpgaPins_Fpga_CPU_is_andi_a3;

// For /fpga_pins/fpga|cpu$is_auipc.
logic FpgaPins_Fpga_CPU_is_auipc_a1,
      FpgaPins_Fpga_CPU_is_auipc_a2,
      FpgaPins_Fpga_CPU_is_auipc_a3;

// For /fpga_pins/fpga|cpu$is_b_instr.
logic FpgaPins_Fpga_CPU_is_b_instr_a1;

// For /fpga_pins/fpga|cpu$is_beq.
logic FpgaPins_Fpga_CPU_is_beq_a1,
      FpgaPins_Fpga_CPU_is_beq_a2,
      FpgaPins_Fpga_CPU_is_beq_a3;

// For /fpga_pins/fpga|cpu$is_bge.
logic FpgaPins_Fpga_CPU_is_bge_a1,
      FpgaPins_Fpga_CPU_is_bge_a2,
      FpgaPins_Fpga_CPU_is_bge_a3;

// For /fpga_pins/fpga|cpu$is_bgeu.
logic FpgaPins_Fpga_CPU_is_bgeu_a1,
      FpgaPins_Fpga_CPU_is_bgeu_a2,
      FpgaPins_Fpga_CPU_is_bgeu_a3;

// For /fpga_pins/fpga|cpu$is_blt.
logic FpgaPins_Fpga_CPU_is_blt_a1,
      FpgaPins_Fpga_CPU_is_blt_a2,
      FpgaPins_Fpga_CPU_is_blt_a3;

// For /fpga_pins/fpga|cpu$is_bltu.
logic FpgaPins_Fpga_CPU_is_bltu_a1,
      FpgaPins_Fpga_CPU_is_bltu_a2,
      FpgaPins_Fpga_CPU_is_bltu_a3;

// For /fpga_pins/fpga|cpu$is_bne.
logic FpgaPins_Fpga_CPU_is_bne_a1,
      FpgaPins_Fpga_CPU_is_bne_a2,
      FpgaPins_Fpga_CPU_is_bne_a3;

// For /fpga_pins/fpga|cpu$is_i_instr.
logic FpgaPins_Fpga_CPU_is_i_instr_a1;

// For /fpga_pins/fpga|cpu$is_j_instr.
logic FpgaPins_Fpga_CPU_is_j_instr_a1;

// For /fpga_pins/fpga|cpu$is_jal.
logic FpgaPins_Fpga_CPU_is_jal_a1,
      FpgaPins_Fpga_CPU_is_jal_a2,
      FpgaPins_Fpga_CPU_is_jal_a3;

// For /fpga_pins/fpga|cpu$is_jalr.
logic FpgaPins_Fpga_CPU_is_jalr_a1,
      FpgaPins_Fpga_CPU_is_jalr_a2,
      FpgaPins_Fpga_CPU_is_jalr_a3;

// For /fpga_pins/fpga|cpu$is_jump.
logic FpgaPins_Fpga_CPU_is_jump_a3;

// For /fpga_pins/fpga|cpu$is_load.
logic FpgaPins_Fpga_CPU_is_load_a1,
      FpgaPins_Fpga_CPU_is_load_a2,
      FpgaPins_Fpga_CPU_is_load_a3,
      FpgaPins_Fpga_CPU_is_load_a4;

// For /fpga_pins/fpga|cpu$is_lui.
logic FpgaPins_Fpga_CPU_is_lui_a1,
      FpgaPins_Fpga_CPU_is_lui_a2,
      FpgaPins_Fpga_CPU_is_lui_a3;

// For /fpga_pins/fpga|cpu$is_or.
logic FpgaPins_Fpga_CPU_is_or_a1,
      FpgaPins_Fpga_CPU_is_or_a2,
      FpgaPins_Fpga_CPU_is_or_a3;

// For /fpga_pins/fpga|cpu$is_ori.
logic FpgaPins_Fpga_CPU_is_ori_a1,
      FpgaPins_Fpga_CPU_is_ori_a2,
      FpgaPins_Fpga_CPU_is_ori_a3;

// For /fpga_pins/fpga|cpu$is_r_instr.
logic FpgaPins_Fpga_CPU_is_r_instr_a1;

// For /fpga_pins/fpga|cpu$is_s_instr.
logic FpgaPins_Fpga_CPU_is_s_instr_a1,
      FpgaPins_Fpga_CPU_is_s_instr_a2,
      FpgaPins_Fpga_CPU_is_s_instr_a3,
      FpgaPins_Fpga_CPU_is_s_instr_a4;

// For /fpga_pins/fpga|cpu$is_sll.
logic FpgaPins_Fpga_CPU_is_sll_a1,
      FpgaPins_Fpga_CPU_is_sll_a2,
      FpgaPins_Fpga_CPU_is_sll_a3;

// For /fpga_pins/fpga|cpu$is_slli.
logic FpgaPins_Fpga_CPU_is_slli_a1,
      FpgaPins_Fpga_CPU_is_slli_a2,
      FpgaPins_Fpga_CPU_is_slli_a3;

// For /fpga_pins/fpga|cpu$is_slt.
logic FpgaPins_Fpga_CPU_is_slt_a1,
      FpgaPins_Fpga_CPU_is_slt_a2,
      FpgaPins_Fpga_CPU_is_slt_a3;

// For /fpga_pins/fpga|cpu$is_slti.
logic FpgaPins_Fpga_CPU_is_slti_a1,
      FpgaPins_Fpga_CPU_is_slti_a2,
      FpgaPins_Fpga_CPU_is_slti_a3;

// For /fpga_pins/fpga|cpu$is_sltiu.
logic FpgaPins_Fpga_CPU_is_sltiu_a1,
      FpgaPins_Fpga_CPU_is_sltiu_a2,
      FpgaPins_Fpga_CPU_is_sltiu_a3;

// For /fpga_pins/fpga|cpu$is_sltu.
logic FpgaPins_Fpga_CPU_is_sltu_a1,
      FpgaPins_Fpga_CPU_is_sltu_a2,
      FpgaPins_Fpga_CPU_is_sltu_a3;

// For /fpga_pins/fpga|cpu$is_sra.
logic FpgaPins_Fpga_CPU_is_sra_a1,
      FpgaPins_Fpga_CPU_is_sra_a2,
      FpgaPins_Fpga_CPU_is_sra_a3;

// For /fpga_pins/fpga|cpu$is_srai.
logic FpgaPins_Fpga_CPU_is_srai_a1,
      FpgaPins_Fpga_CPU_is_srai_a2,
      FpgaPins_Fpga_CPU_is_srai_a3;

// For /fpga_pins/fpga|cpu$is_srl.
logic FpgaPins_Fpga_CPU_is_srl_a1,
      FpgaPins_Fpga_CPU_is_srl_a2,
      FpgaPins_Fpga_CPU_is_srl_a3;

// For /fpga_pins/fpga|cpu$is_srli.
logic FpgaPins_Fpga_CPU_is_srli_a1,
      FpgaPins_Fpga_CPU_is_srli_a2,
      FpgaPins_Fpga_CPU_is_srli_a3;

// For /fpga_pins/fpga|cpu$is_sub.
logic FpgaPins_Fpga_CPU_is_sub_a1,
      FpgaPins_Fpga_CPU_is_sub_a2,
      FpgaPins_Fpga_CPU_is_sub_a3;

// For /fpga_pins/fpga|cpu$is_u_instr.
logic FpgaPins_Fpga_CPU_is_u_instr_a1;

// For /fpga_pins/fpga|cpu$is_xor.
logic FpgaPins_Fpga_CPU_is_xor_a1,
      FpgaPins_Fpga_CPU_is_xor_a2,
      FpgaPins_Fpga_CPU_is_xor_a3;

// For /fpga_pins/fpga|cpu$is_xori.
logic FpgaPins_Fpga_CPU_is_xori_a1,
      FpgaPins_Fpga_CPU_is_xori_a2,
      FpgaPins_Fpga_CPU_is_xori_a3;

// For /fpga_pins/fpga|cpu$jalr_tgt_pc.
logic [31:0] FpgaPins_Fpga_CPU_jalr_tgt_pc_a3;

// For /fpga_pins/fpga|cpu$ld_data.
logic [31:0] FpgaPins_Fpga_CPU_ld_data_a5;

// For /fpga_pins/fpga|cpu$opcode.
logic [6:0] FpgaPins_Fpga_CPU_opcode_a1;

// For /fpga_pins/fpga|cpu$pc.
logic [31:0] FpgaPins_Fpga_CPU_pc_a0,
             FpgaPins_Fpga_CPU_pc_a1,
             FpgaPins_Fpga_CPU_pc_a2,
             FpgaPins_Fpga_CPU_pc_a3;

// For /fpga_pins/fpga|cpu$rd.
logic [4:0] FpgaPins_Fpga_CPU_rd_a1,
            FpgaPins_Fpga_CPU_rd_a2,
            FpgaPins_Fpga_CPU_rd_a3,
            FpgaPins_Fpga_CPU_rd_a4,
            FpgaPins_Fpga_CPU_rd_a5;

// For /fpga_pins/fpga|cpu$rd_valid.
logic FpgaPins_Fpga_CPU_rd_valid_a1,
      FpgaPins_Fpga_CPU_rd_valid_a2,
      FpgaPins_Fpga_CPU_rd_valid_a3;

// For /fpga_pins/fpga|cpu$reset.
logic FpgaPins_Fpga_CPU_reset_a0,
      FpgaPins_Fpga_CPU_reset_a1,
      FpgaPins_Fpga_CPU_reset_a2,
      FpgaPins_Fpga_CPU_reset_a3,
      FpgaPins_Fpga_CPU_reset_a4;

// For /fpga_pins/fpga|cpu$result.
logic [31:0] FpgaPins_Fpga_CPU_result_a3;
logic [4:2] FpgaPins_Fpga_CPU_result_a4;

// For /fpga_pins/fpga|cpu$rf_rd_data1.
logic [31:0] FpgaPins_Fpga_CPU_rf_rd_data1_a2;

// For /fpga_pins/fpga|cpu$rf_rd_data2.
logic [31:0] FpgaPins_Fpga_CPU_rf_rd_data2_a2;

// For /fpga_pins/fpga|cpu$rf_rd_en1.
logic FpgaPins_Fpga_CPU_rf_rd_en1_a2;

// For /fpga_pins/fpga|cpu$rf_rd_en2.
logic FpgaPins_Fpga_CPU_rf_rd_en2_a2;

// For /fpga_pins/fpga|cpu$rf_rd_index1.
logic [4:0] FpgaPins_Fpga_CPU_rf_rd_index1_a2;

// For /fpga_pins/fpga|cpu$rf_rd_index2.
logic [4:0] FpgaPins_Fpga_CPU_rf_rd_index2_a2;

// For /fpga_pins/fpga|cpu$rf_wr_data.
logic [31:0] FpgaPins_Fpga_CPU_rf_wr_data_a3;

// For /fpga_pins/fpga|cpu$rf_wr_en.
logic FpgaPins_Fpga_CPU_rf_wr_en_a3;

// For /fpga_pins/fpga|cpu$rf_wr_index.
logic [4:0] FpgaPins_Fpga_CPU_rf_wr_index_a3;

// For /fpga_pins/fpga|cpu$rs1.
logic [4:0] FpgaPins_Fpga_CPU_rs1_a1,
            FpgaPins_Fpga_CPU_rs1_a2;

// For /fpga_pins/fpga|cpu$rs1_valid.
logic FpgaPins_Fpga_CPU_rs1_valid_a1,
      FpgaPins_Fpga_CPU_rs1_valid_a2;

// For /fpga_pins/fpga|cpu$rs2.
logic [4:0] FpgaPins_Fpga_CPU_rs2_a1,
            FpgaPins_Fpga_CPU_rs2_a2;

// For /fpga_pins/fpga|cpu$rs2_valid.
logic FpgaPins_Fpga_CPU_rs2_valid_a1,
      FpgaPins_Fpga_CPU_rs2_valid_a2;

// For /fpga_pins/fpga|cpu$sltiu_rslt.
logic [31:0] FpgaPins_Fpga_CPU_sltiu_rslt_a3;

// For /fpga_pins/fpga|cpu$sltu_rslt.
logic [31:0] FpgaPins_Fpga_CPU_sltu_rslt_a3;

// For /fpga_pins/fpga|cpu$src1_value.
logic [31:0] FpgaPins_Fpga_CPU_src1_value_a2,
             FpgaPins_Fpga_CPU_src1_value_a3;

// For /fpga_pins/fpga|cpu$src2_value.
logic [31:0] FpgaPins_Fpga_CPU_src2_value_a2,
             FpgaPins_Fpga_CPU_src2_value_a3,
             FpgaPins_Fpga_CPU_src2_value_a4;

// For /fpga_pins/fpga|cpu$taken_br.
logic FpgaPins_Fpga_CPU_taken_br_a3;

// For /fpga_pins/fpga|cpu$valid.
logic FpgaPins_Fpga_CPU_valid_a3,
      FpgaPins_Fpga_CPU_valid_a4;

// For /fpga_pins/fpga|cpu$valid_jump.
logic FpgaPins_Fpga_CPU_valid_jump_a3,
      FpgaPins_Fpga_CPU_valid_jump_a4,
      FpgaPins_Fpga_CPU_valid_jump_a5;

// For /fpga_pins/fpga|cpu$valid_load.
logic FpgaPins_Fpga_CPU_valid_load_a3,
      FpgaPins_Fpga_CPU_valid_load_a4,
      FpgaPins_Fpga_CPU_valid_load_a5;

// For /fpga_pins/fpga|cpu$valid_taken_br.
logic FpgaPins_Fpga_CPU_valid_taken_br_a3,
      FpgaPins_Fpga_CPU_valid_taken_br_a4,
      FpgaPins_Fpga_CPU_valid_taken_br_a5;

// For /fpga_pins/fpga|cpu/dmem$value.
logic [31:0] FpgaPins_Fpga_CPU_Dmem_value_a4 [7:0],
             FpgaPins_Fpga_CPU_Dmem_value_a5 [7:0];

// For /fpga_pins/fpga|cpu/imem$instr.
logic [31:0] FpgaPins_Fpga_CPU_Imem_instr_a1 [9:0];

// For /fpga_pins/fpga|cpu/xreg$value.
logic [31:0] FpgaPins_Fpga_CPU_Xreg_value_a3 [15:0],
             FpgaPins_Fpga_CPU_Xreg_value_a4 [15:0],
             FpgaPins_Fpga_CPU_Xreg_value_a5 [15:0],
             FpgaPins_Fpga_CPU_Xreg_value_a6 [15:0];




   //
   // Scope: /fpga_pins
   //


      //
      // Scope: /fpga
      //


         //
         // Scope: |cpu
         //

            // Staging of $br_tgt_pc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_br_tgt_pc_a3[31:0] <= FpgaPins_Fpga_CPU_br_tgt_pc_a2[31:0];

            // Staging of $dmem_rd_data.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_dmem_rd_data_a5[31:0] <= FpgaPins_Fpga_CPU_dmem_rd_data_a4[31:0];

            // Staging of $imem_rd_addr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_imem_rd_addr_a1[4-1:0] <= FpgaPins_Fpga_CPU_imem_rd_addr_a0[4-1:0];

            // Staging of $imem_rd_en.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_imem_rd_en_a1 <= FpgaPins_Fpga_CPU_imem_rd_en_a0;

            // Staging of $imm.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_imm_a2[31:0] <= FpgaPins_Fpga_CPU_imm_a1[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_imm_a3[31:0] <= FpgaPins_Fpga_CPU_imm_a2[31:0];

            // Staging of $inc_pc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_inc_pc_a2[31:0] <= FpgaPins_Fpga_CPU_inc_pc_a1[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_inc_pc_a3[31:0] <= FpgaPins_Fpga_CPU_inc_pc_a2[31:0];

            // Staging of $is_add.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_add_a2 <= FpgaPins_Fpga_CPU_is_add_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_add_a3 <= FpgaPins_Fpga_CPU_is_add_a2;

            // Staging of $is_addi.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_addi_a2 <= FpgaPins_Fpga_CPU_is_addi_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_addi_a3 <= FpgaPins_Fpga_CPU_is_addi_a2;

            // Staging of $is_and.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_and_a2 <= FpgaPins_Fpga_CPU_is_and_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_and_a3 <= FpgaPins_Fpga_CPU_is_and_a2;

            // Staging of $is_andi.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_andi_a2 <= FpgaPins_Fpga_CPU_is_andi_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_andi_a3 <= FpgaPins_Fpga_CPU_is_andi_a2;

            // Staging of $is_auipc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_auipc_a2 <= FpgaPins_Fpga_CPU_is_auipc_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_auipc_a3 <= FpgaPins_Fpga_CPU_is_auipc_a2;

            // Staging of $is_beq.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_beq_a2 <= FpgaPins_Fpga_CPU_is_beq_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_beq_a3 <= FpgaPins_Fpga_CPU_is_beq_a2;

            // Staging of $is_bge.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bge_a2 <= FpgaPins_Fpga_CPU_is_bge_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bge_a3 <= FpgaPins_Fpga_CPU_is_bge_a2;

            // Staging of $is_bgeu.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bgeu_a2 <= FpgaPins_Fpga_CPU_is_bgeu_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bgeu_a3 <= FpgaPins_Fpga_CPU_is_bgeu_a2;

            // Staging of $is_blt.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_blt_a2 <= FpgaPins_Fpga_CPU_is_blt_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_blt_a3 <= FpgaPins_Fpga_CPU_is_blt_a2;

            // Staging of $is_bltu.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bltu_a2 <= FpgaPins_Fpga_CPU_is_bltu_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bltu_a3 <= FpgaPins_Fpga_CPU_is_bltu_a2;

            // Staging of $is_bne.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bne_a2 <= FpgaPins_Fpga_CPU_is_bne_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_bne_a3 <= FpgaPins_Fpga_CPU_is_bne_a2;

            // Staging of $is_jal.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jal_a2 <= FpgaPins_Fpga_CPU_is_jal_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jal_a3 <= FpgaPins_Fpga_CPU_is_jal_a2;

            // Staging of $is_jalr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jalr_a2 <= FpgaPins_Fpga_CPU_is_jalr_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_jalr_a3 <= FpgaPins_Fpga_CPU_is_jalr_a2;

            // Staging of $is_load.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_load_a2 <= FpgaPins_Fpga_CPU_is_load_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_load_a3 <= FpgaPins_Fpga_CPU_is_load_a2;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_load_a4 <= FpgaPins_Fpga_CPU_is_load_a3;

            // Staging of $is_lui.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_lui_a2 <= FpgaPins_Fpga_CPU_is_lui_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_lui_a3 <= FpgaPins_Fpga_CPU_is_lui_a2;

            // Staging of $is_or.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_or_a2 <= FpgaPins_Fpga_CPU_is_or_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_or_a3 <= FpgaPins_Fpga_CPU_is_or_a2;

            // Staging of $is_ori.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_ori_a2 <= FpgaPins_Fpga_CPU_is_ori_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_ori_a3 <= FpgaPins_Fpga_CPU_is_ori_a2;

            // Staging of $is_s_instr.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_s_instr_a2 <= FpgaPins_Fpga_CPU_is_s_instr_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_s_instr_a3 <= FpgaPins_Fpga_CPU_is_s_instr_a2;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_s_instr_a4 <= FpgaPins_Fpga_CPU_is_s_instr_a3;

            // Staging of $is_sll.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sll_a2 <= FpgaPins_Fpga_CPU_is_sll_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sll_a3 <= FpgaPins_Fpga_CPU_is_sll_a2;

            // Staging of $is_slli.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slli_a2 <= FpgaPins_Fpga_CPU_is_slli_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slli_a3 <= FpgaPins_Fpga_CPU_is_slli_a2;

            // Staging of $is_slt.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slt_a2 <= FpgaPins_Fpga_CPU_is_slt_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slt_a3 <= FpgaPins_Fpga_CPU_is_slt_a2;

            // Staging of $is_slti.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slti_a2 <= FpgaPins_Fpga_CPU_is_slti_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_slti_a3 <= FpgaPins_Fpga_CPU_is_slti_a2;

            // Staging of $is_sltiu.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sltiu_a2 <= FpgaPins_Fpga_CPU_is_sltiu_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sltiu_a3 <= FpgaPins_Fpga_CPU_is_sltiu_a2;

            // Staging of $is_sltu.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sltu_a2 <= FpgaPins_Fpga_CPU_is_sltu_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sltu_a3 <= FpgaPins_Fpga_CPU_is_sltu_a2;

            // Staging of $is_sra.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sra_a2 <= FpgaPins_Fpga_CPU_is_sra_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sra_a3 <= FpgaPins_Fpga_CPU_is_sra_a2;

            // Staging of $is_srai.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srai_a2 <= FpgaPins_Fpga_CPU_is_srai_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srai_a3 <= FpgaPins_Fpga_CPU_is_srai_a2;

            // Staging of $is_srl.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srl_a2 <= FpgaPins_Fpga_CPU_is_srl_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srl_a3 <= FpgaPins_Fpga_CPU_is_srl_a2;

            // Staging of $is_srli.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srli_a2 <= FpgaPins_Fpga_CPU_is_srli_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_srli_a3 <= FpgaPins_Fpga_CPU_is_srli_a2;

            // Staging of $is_sub.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sub_a2 <= FpgaPins_Fpga_CPU_is_sub_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_sub_a3 <= FpgaPins_Fpga_CPU_is_sub_a2;

            // Staging of $is_xor.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_xor_a2 <= FpgaPins_Fpga_CPU_is_xor_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_xor_a3 <= FpgaPins_Fpga_CPU_is_xor_a2;

            // Staging of $is_xori.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_xori_a2 <= FpgaPins_Fpga_CPU_is_xori_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_is_xori_a3 <= FpgaPins_Fpga_CPU_is_xori_a2;

            // Staging of $pc.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_pc_a1[31:0] <= FpgaPins_Fpga_CPU_pc_a0[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_pc_a2[31:0] <= FpgaPins_Fpga_CPU_pc_a1[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_pc_a3[31:0] <= FpgaPins_Fpga_CPU_pc_a2[31:0];

            // Staging of $rd.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a2[4:0] <= FpgaPins_Fpga_CPU_rd_a1[4:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a3[4:0] <= FpgaPins_Fpga_CPU_rd_a2[4:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a4[4:0] <= FpgaPins_Fpga_CPU_rd_a3[4:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_a5[4:0] <= FpgaPins_Fpga_CPU_rd_a4[4:0];

            // Staging of $rd_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_valid_a2 <= FpgaPins_Fpga_CPU_rd_valid_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rd_valid_a3 <= FpgaPins_Fpga_CPU_rd_valid_a2;

            // Staging of $reset.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a1 <= FpgaPins_Fpga_CPU_reset_a0;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a2 <= FpgaPins_Fpga_CPU_reset_a1;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a3 <= FpgaPins_Fpga_CPU_reset_a2;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_reset_a4 <= FpgaPins_Fpga_CPU_reset_a3;

            // Staging of $result.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_result_a4[4:2] <= FpgaPins_Fpga_CPU_result_a3[4:2];

            // Staging of $rs1.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs1_a2[4:0] <= FpgaPins_Fpga_CPU_rs1_a1[4:0];

            // Staging of $rs1_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs1_valid_a2 <= FpgaPins_Fpga_CPU_rs1_valid_a1;

            // Staging of $rs2.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs2_a2[4:0] <= FpgaPins_Fpga_CPU_rs2_a1[4:0];

            // Staging of $rs2_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_rs2_valid_a2 <= FpgaPins_Fpga_CPU_rs2_valid_a1;

            // Staging of $src1_value.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_src1_value_a3[31:0] <= FpgaPins_Fpga_CPU_src1_value_a2[31:0];

            // Staging of $src2_value.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_src2_value_a3[31:0] <= FpgaPins_Fpga_CPU_src2_value_a2[31:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_src2_value_a4[31:0] <= FpgaPins_Fpga_CPU_src2_value_a3[31:0];

            // Staging of $valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_a4 <= FpgaPins_Fpga_CPU_valid_a3;

            // Staging of $valid_jump.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_jump_a4 <= FpgaPins_Fpga_CPU_valid_jump_a3;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_jump_a5 <= FpgaPins_Fpga_CPU_valid_jump_a4;

            // Staging of $valid_load.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_load_a4 <= FpgaPins_Fpga_CPU_valid_load_a3;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_load_a5 <= FpgaPins_Fpga_CPU_valid_load_a4;

            // Staging of $valid_taken_br.
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_taken_br_a4 <= FpgaPins_Fpga_CPU_valid_taken_br_a3;
            always_ff @(posedge clk) FpgaPins_Fpga_CPU_valid_taken_br_a5 <= FpgaPins_Fpga_CPU_valid_taken_br_a4;


            //
            // Scope: /dmem[7:0]
            //
            for (dmem = 0; dmem <= 7; dmem++) begin : L1gen_FpgaPins_Fpga_CPU_Dmem
               // Staging of $value.
               always_ff @(posedge clk) FpgaPins_Fpga_CPU_Dmem_value_a5[dmem][31:0] <= FpgaPins_Fpga_CPU_Dmem_value_a4[dmem][31:0];

            end

            //
            // Scope: /xreg[15:0]
            //
            for (xreg = 0; xreg <= 15; xreg++) begin : L1gen_FpgaPins_Fpga_CPU_Xreg
               // Staging of $value.
               always_ff @(posedge clk) FpgaPins_Fpga_CPU_Xreg_value_a4[xreg][31:0] <= FpgaPins_Fpga_CPU_Xreg_value_a3[xreg][31:0];
               always_ff @(posedge clk) FpgaPins_Fpga_CPU_Xreg_value_a5[xreg][31:0] <= FpgaPins_Fpga_CPU_Xreg_value_a4[xreg][31:0];
               always_ff @(posedge clk) FpgaPins_Fpga_CPU_Xreg_value_a6[xreg][31:0] <= FpgaPins_Fpga_CPU_Xreg_value_a5[xreg][31:0];

            end







//
// Debug Signals
//

   if (1) begin : DEBUG_SIGS_GTKWAVE

      (* keep *) logic [7:0] \@0$slideswitch ;
      assign \@0$slideswitch = L0_slideswitch_a0;
      (* keep *) logic  \@0$sseg_decimal_point_n ;
      assign \@0$sseg_decimal_point_n = L0_sseg_decimal_point_n_a0;
      (* keep *) logic [7:0] \@0$sseg_digit_n ;
      assign \@0$sseg_digit_n = L0_sseg_digit_n_a0;
      (* keep *) logic [6:0] \@0$sseg_segment_n ;
      assign \@0$sseg_segment_n = L0_sseg_segment_n_a0;

      //
      // Scope: /digit[0:0]
      //
      for (digit = 0; digit <= 0; digit++) begin : \/digit 

         //
         // Scope: /leds[7:0]
         //
         for (leds = 0; leds <= 7; leds++) begin : \/leds 
            (* keep *) logic  \//@0$viz_lit ;
            assign \//@0$viz_lit = L1_Digit[digit].L2_Leds[leds].L2_viz_lit_a0;
         end
      end

      //
      // Scope: /fpga_pins
      //
      if (1) begin : \/fpga_pins 

         //
         // Scope: /fpga
         //
         if (1) begin : \/fpga 

            //
            // Scope: |cpu
            //
            if (1) begin : P_cpu
               (* keep *) logic [31:0] \///@2$br_tgt_pc ;
               assign \///@2$br_tgt_pc = FpgaPins_Fpga_CPU_br_tgt_pc_a2;
               (* keep *) logic [10:0] \///@1$dec_bits ;
               assign \///@1$dec_bits = FpgaPins_Fpga_CPU_dec_bits_a1;
               (* keep *) logic [2:0] \///@4$dmem_addr ;
               assign \///@4$dmem_addr = FpgaPins_Fpga_CPU_dmem_addr_a4;
               (* keep *) logic [31:0] \///?$dmem_rd_en@4$dmem_rd_data ;
               assign \///?$dmem_rd_en@4$dmem_rd_data = FpgaPins_Fpga_CPU_dmem_rd_data_a4;
               (* keep *) logic  \///@4$dmem_rd_en ;
               assign \///@4$dmem_rd_en = FpgaPins_Fpga_CPU_dmem_rd_en_a4;
               (* keep *) logic [31:0] \///@4$dmem_wr_data ;
               assign \///@4$dmem_wr_data = FpgaPins_Fpga_CPU_dmem_wr_data_a4;
               (* keep *) logic  \///@4$dmem_wr_en ;
               assign \///@4$dmem_wr_en = FpgaPins_Fpga_CPU_dmem_wr_en_a4;
               (* keep *) logic [2:0] \///?$funct3_valid@1$funct3 ;
               assign \///?$funct3_valid@1$funct3 = FpgaPins_Fpga_CPU_funct3_a1;
               (* keep *) logic  \///@1$funct3_valid ;
               assign \///@1$funct3_valid = FpgaPins_Fpga_CPU_funct3_valid_a1;
               (* keep *) logic [6:0] \///?$funct7_valid@1$funct7 ;
               assign \///?$funct7_valid@1$funct7 = FpgaPins_Fpga_CPU_funct7_a1;
               (* keep *) logic  \///@1$funct7_valid ;
               assign \///@1$funct7_valid = FpgaPins_Fpga_CPU_funct7_valid_a1;
               (* keep *) logic [4-1:0] \///@0$imem_rd_addr ;
               assign \///@0$imem_rd_addr = FpgaPins_Fpga_CPU_imem_rd_addr_a0;
               (* keep *) logic [31:0] \///?$imem_rd_en@1$imem_rd_data ;
               assign \///?$imem_rd_en@1$imem_rd_data = FpgaPins_Fpga_CPU_imem_rd_data_a1;
               (* keep *) logic  \///@0$imem_rd_en ;
               assign \///@0$imem_rd_en = FpgaPins_Fpga_CPU_imem_rd_en_a0;
               (* keep *) logic [31:0] \///@1$imm ;
               assign \///@1$imm = FpgaPins_Fpga_CPU_imm_a1;
               (* keep *) logic [31:0] \///@1$inc_pc ;
               assign \///@1$inc_pc = FpgaPins_Fpga_CPU_inc_pc_a1;
               (* keep *) logic [31:0] \///@1$instr ;
               assign \///@1$instr = FpgaPins_Fpga_CPU_instr_a1;
               (* keep *) logic  \///@1$is_add ;
               assign \///@1$is_add = FpgaPins_Fpga_CPU_is_add_a1;
               (* keep *) logic  \///@1$is_addi ;
               assign \///@1$is_addi = FpgaPins_Fpga_CPU_is_addi_a1;
               (* keep *) logic  \///@1$is_and ;
               assign \///@1$is_and = FpgaPins_Fpga_CPU_is_and_a1;
               (* keep *) logic  \///@1$is_andi ;
               assign \///@1$is_andi = FpgaPins_Fpga_CPU_is_andi_a1;
               (* keep *) logic  \///@1$is_auipc ;
               assign \///@1$is_auipc = FpgaPins_Fpga_CPU_is_auipc_a1;
               (* keep *) logic  \///@1$is_b_instr ;
               assign \///@1$is_b_instr = FpgaPins_Fpga_CPU_is_b_instr_a1;
               (* keep *) logic  \///@1$is_beq ;
               assign \///@1$is_beq = FpgaPins_Fpga_CPU_is_beq_a1;
               (* keep *) logic  \///@1$is_bge ;
               assign \///@1$is_bge = FpgaPins_Fpga_CPU_is_bge_a1;
               (* keep *) logic  \///@1$is_bgeu ;
               assign \///@1$is_bgeu = FpgaPins_Fpga_CPU_is_bgeu_a1;
               (* keep *) logic  \///@1$is_blt ;
               assign \///@1$is_blt = FpgaPins_Fpga_CPU_is_blt_a1;
               (* keep *) logic  \///@1$is_bltu ;
               assign \///@1$is_bltu = FpgaPins_Fpga_CPU_is_bltu_a1;
               (* keep *) logic  \///@1$is_bne ;
               assign \///@1$is_bne = FpgaPins_Fpga_CPU_is_bne_a1;
               (* keep *) logic  \///@1$is_i_instr ;
               assign \///@1$is_i_instr = FpgaPins_Fpga_CPU_is_i_instr_a1;
               (* keep *) logic  \///@1$is_j_instr ;
               assign \///@1$is_j_instr = FpgaPins_Fpga_CPU_is_j_instr_a1;
               (* keep *) logic  \///@1$is_jal ;
               assign \///@1$is_jal = FpgaPins_Fpga_CPU_is_jal_a1;
               (* keep *) logic  \///@1$is_jalr ;
               assign \///@1$is_jalr = FpgaPins_Fpga_CPU_is_jalr_a1;
               (* keep *) logic  \///@3$is_jump ;
               assign \///@3$is_jump = FpgaPins_Fpga_CPU_is_jump_a3;
               (* keep *) logic  \///@1$is_load ;
               assign \///@1$is_load = FpgaPins_Fpga_CPU_is_load_a1;
               (* keep *) logic  \///@1$is_lui ;
               assign \///@1$is_lui = FpgaPins_Fpga_CPU_is_lui_a1;
               (* keep *) logic  \///@1$is_or ;
               assign \///@1$is_or = FpgaPins_Fpga_CPU_is_or_a1;
               (* keep *) logic  \///@1$is_ori ;
               assign \///@1$is_ori = FpgaPins_Fpga_CPU_is_ori_a1;
               (* keep *) logic  \///@1$is_r_instr ;
               assign \///@1$is_r_instr = FpgaPins_Fpga_CPU_is_r_instr_a1;
               (* keep *) logic  \///@1$is_s_instr ;
               assign \///@1$is_s_instr = FpgaPins_Fpga_CPU_is_s_instr_a1;
               (* keep *) logic  \///@1$is_sll ;
               assign \///@1$is_sll = FpgaPins_Fpga_CPU_is_sll_a1;
               (* keep *) logic  \///@1$is_slli ;
               assign \///@1$is_slli = FpgaPins_Fpga_CPU_is_slli_a1;
               (* keep *) logic  \///@1$is_slt ;
               assign \///@1$is_slt = FpgaPins_Fpga_CPU_is_slt_a1;
               (* keep *) logic  \///@1$is_slti ;
               assign \///@1$is_slti = FpgaPins_Fpga_CPU_is_slti_a1;
               (* keep *) logic  \///@1$is_sltiu ;
               assign \///@1$is_sltiu = FpgaPins_Fpga_CPU_is_sltiu_a1;
               (* keep *) logic  \///@1$is_sltu ;
               assign \///@1$is_sltu = FpgaPins_Fpga_CPU_is_sltu_a1;
               (* keep *) logic  \///@1$is_sra ;
               assign \///@1$is_sra = FpgaPins_Fpga_CPU_is_sra_a1;
               (* keep *) logic  \///@1$is_srai ;
               assign \///@1$is_srai = FpgaPins_Fpga_CPU_is_srai_a1;
               (* keep *) logic  \///@1$is_srl ;
               assign \///@1$is_srl = FpgaPins_Fpga_CPU_is_srl_a1;
               (* keep *) logic  \///@1$is_srli ;
               assign \///@1$is_srli = FpgaPins_Fpga_CPU_is_srli_a1;
               (* keep *) logic  \///@1$is_sub ;
               assign \///@1$is_sub = FpgaPins_Fpga_CPU_is_sub_a1;
               (* keep *) logic  \///@1$is_u_instr ;
               assign \///@1$is_u_instr = FpgaPins_Fpga_CPU_is_u_instr_a1;
               (* keep *) logic  \///@1$is_xor ;
               assign \///@1$is_xor = FpgaPins_Fpga_CPU_is_xor_a1;
               (* keep *) logic  \///@1$is_xori ;
               assign \///@1$is_xori = FpgaPins_Fpga_CPU_is_xori_a1;
               (* keep *) logic [31:0] \///@3$jalr_tgt_pc ;
               assign \///@3$jalr_tgt_pc = FpgaPins_Fpga_CPU_jalr_tgt_pc_a3;
               (* keep *) logic [31:0] \///@5$ld_data ;
               assign \///@5$ld_data = FpgaPins_Fpga_CPU_ld_data_a5;
               (* keep *) logic [6:0] \///@1$opcode ;
               assign \///@1$opcode = FpgaPins_Fpga_CPU_opcode_a1;
               (* keep *) logic [31:0] \///@0$pc ;
               assign \///@0$pc = FpgaPins_Fpga_CPU_pc_a0;
               (* keep *) logic [4:0] \///?$rd_valid@1$rd ;
               assign \///?$rd_valid@1$rd = FpgaPins_Fpga_CPU_rd_a1;
               (* keep *) logic  \///@1$rd_valid ;
               assign \///@1$rd_valid = FpgaPins_Fpga_CPU_rd_valid_a1;
               (* keep *) logic  \///@0$reset ;
               assign \///@0$reset = FpgaPins_Fpga_CPU_reset_a0;
               (* keep *) logic [31:0] \///@3$result ;
               assign \///@3$result = FpgaPins_Fpga_CPU_result_a3;
               (* keep *) logic [31:0] \///?$rf_rd_en1@2$rf_rd_data1 ;
               assign \///?$rf_rd_en1@2$rf_rd_data1 = FpgaPins_Fpga_CPU_rf_rd_data1_a2;
               (* keep *) logic [31:0] \///?$rf_rd_en2@2$rf_rd_data2 ;
               assign \///?$rf_rd_en2@2$rf_rd_data2 = FpgaPins_Fpga_CPU_rf_rd_data2_a2;
               (* keep *) logic  \///@2$rf_rd_en1 ;
               assign \///@2$rf_rd_en1 = FpgaPins_Fpga_CPU_rf_rd_en1_a2;
               (* keep *) logic  \///@2$rf_rd_en2 ;
               assign \///@2$rf_rd_en2 = FpgaPins_Fpga_CPU_rf_rd_en2_a2;
               (* keep *) logic [4:0] \///@2$rf_rd_index1 ;
               assign \///@2$rf_rd_index1 = FpgaPins_Fpga_CPU_rf_rd_index1_a2;
               (* keep *) logic [4:0] \///@2$rf_rd_index2 ;
               assign \///@2$rf_rd_index2 = FpgaPins_Fpga_CPU_rf_rd_index2_a2;
               (* keep *) logic [31:0] \///@3$rf_wr_data ;
               assign \///@3$rf_wr_data = FpgaPins_Fpga_CPU_rf_wr_data_a3;
               (* keep *) logic  \///@3$rf_wr_en ;
               assign \///@3$rf_wr_en = FpgaPins_Fpga_CPU_rf_wr_en_a3;
               (* keep *) logic [4:0] \///@3$rf_wr_index ;
               assign \///@3$rf_wr_index = FpgaPins_Fpga_CPU_rf_wr_index_a3;
               (* keep *) logic [4:0] \///?$rs1_valid@1$rs1 ;
               assign \///?$rs1_valid@1$rs1 = FpgaPins_Fpga_CPU_rs1_a1;
               (* keep *) logic  \///@1$rs1_valid ;
               assign \///@1$rs1_valid = FpgaPins_Fpga_CPU_rs1_valid_a1;
               (* keep *) logic [4:0] \///?$rs2_valid@1$rs2 ;
               assign \///?$rs2_valid@1$rs2 = FpgaPins_Fpga_CPU_rs2_a1;
               (* keep *) logic  \///@1$rs2_valid ;
               assign \///@1$rs2_valid = FpgaPins_Fpga_CPU_rs2_valid_a1;
               (* keep *) logic [31:0] \///@3$sltiu_rslt ;
               assign \///@3$sltiu_rslt = FpgaPins_Fpga_CPU_sltiu_rslt_a3;
               (* keep *) logic [31:0] \///@3$sltu_rslt ;
               assign \///@3$sltu_rslt = FpgaPins_Fpga_CPU_sltu_rslt_a3;
               (* keep *) logic [31:0] \///@2$src1_value ;
               assign \///@2$src1_value = FpgaPins_Fpga_CPU_src1_value_a2;
               (* keep *) logic [31:0] \///@2$src2_value ;
               assign \///@2$src2_value = FpgaPins_Fpga_CPU_src2_value_a2;
               (* keep *) logic  \///@3$taken_br ;
               assign \///@3$taken_br = FpgaPins_Fpga_CPU_taken_br_a3;
               (* keep *) logic  \///@3$valid ;
               assign \///@3$valid = FpgaPins_Fpga_CPU_valid_a3;
               (* keep *) logic  \///@3$valid_jump ;
               assign \///@3$valid_jump = FpgaPins_Fpga_CPU_valid_jump_a3;
               (* keep *) logic  \///@3$valid_load ;
               assign \///@3$valid_load = FpgaPins_Fpga_CPU_valid_load_a3;
               (* keep *) logic  \///@3$valid_taken_br ;
               assign \///@3$valid_taken_br = FpgaPins_Fpga_CPU_valid_taken_br_a3;

               //
               // Scope: /dmem[7:0]
               //
               for (dmem = 0; dmem <= 7; dmem++) begin : \/dmem 
                  (* keep *) logic [31:0] \////@4$value ;
                  assign \////@4$value = FpgaPins_Fpga_CPU_Dmem_value_a4[dmem];
                  (* keep *) logic  \////@4$wr ;
                  assign \////@4$wr = L1_FpgaPins_Fpga_CPU_Dmem[dmem].L1_wr_a4;
               end

               //
               // Scope: /imem[9:0]
               //
               for (imem = 0; imem <= 9; imem++) begin : \/imem 
                  (* keep *) logic [31:0] \////@1$instr ;
                  assign \////@1$instr = FpgaPins_Fpga_CPU_Imem_instr_a1[imem];
               end

               //
               // Scope: /xreg[15:0]
               //
               for (xreg = 0; xreg <= 15; xreg++) begin : \/xreg 
                  (* keep *) logic [31:0] \////@3$value ;
                  assign \////@3$value = FpgaPins_Fpga_CPU_Xreg_value_a3[xreg];
                  (* keep *) logic  \////@3$wr ;
                  assign \////@3$wr = L1_FpgaPins_Fpga_CPU_Xreg[xreg].L1_wr_a3;
               end
            end
         end
      end

      //
      // Scope: /switch[7:0]
      //
      for (switch = 0; switch <= 7; switch++) begin : \/switch 
         (* keep *) logic  \/@0$viz_switch ;
         assign \/@0$viz_switch = L1_Switch[switch].L1_viz_switch_a0;
      end


   end

// ---------- Generated Code Ends ----------
//_\TLV
   /* verilator lint_off UNOPTFLAT */
   // Connect Tiny Tapeout I/Os to Virtual FPGA Lab.
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/af18805ea79802b83477cf86aff503e97ed7394a/tlvlib/tinytapeoutlib.tlv 67   // Instantiated from top.tlv, 858 as: m5+tt_connections()
      assign L0_slideswitch_a0[7:0] = ui_in;
      assign L0_sseg_segment_n_a0[6:0] = uo_out[6:0];
      assign L0_sseg_decimal_point_n_a0 = uo_out[7];
      assign L0_sseg_digit_n_a0[7:0] = 8'b11111110;
   //_\end_source

   // Instantiate the Virtual FPGA Lab.
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 307   // Instantiated from top.tlv, 861 as: m5+board(/top, /fpga, 7, $, , hidden_solution)
      
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 355   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 309 as: m4+thanks(m5__l(309)m5_eval(m5_get(BOARD_THANKS_ARGS)))
         //_/thanks
            
      //_\end_source
      
   
      // Board VIZ.
   
      // Board Image.
      
      //_/fpga_pins
         
         //_/fpga
            //_\source top.tlv 173   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 340 as: m4+hidden_solution.
               //_\source top.tlv 278   // Instantiated from top.tlv, 174 as: m5+call(m5__l(174)m5_call(if,m5_get(CalcLab), calc_solution, cpu_solution))
                  //_\source M5-FN-riscv_gen 0   // Instantiated from top.tlv, 279 as: m5+riscv_gen()
                     
                  //_\end_source
                  //_\source M5-FN-riscv_sum_prog 0   // Instantiated from top.tlv, 280 as: m5+riscv_sum_prog()
                     // Inst #0: ADD x10, x0, x0
                     // Inst #1: ADD x14, x10, x0
                     // Inst #2: ADDI x12, x10, 10
                     // Inst #3: ADD x13, x10, x0
                     // Inst #4: ADD x14, x13, x14
                     // Inst #5: ADDI x13, x13, 1
                     // Inst #6: BLT x13, x12, loop
                     // Inst #7: ADD x10, x14, x0
                     // Inst #8: SW x0, x10, 4
                     // Inst #9: LW x15, x0, 4
                     
                  //_\end_source
                  
                  //_|cpu
                     //_@0
                        assign FpgaPins_Fpga_CPU_reset_a0 = reset;
               
               
                     // ============================================================================================================
                     // Solutions: Cut this section to provide the shell.
               
                     
                     
               
               
                     // Define the logic that will be included, based on lab ID.
                     // Lab m5_get(LabId): Next PC
                     
                     
                     
                     // Lab m5_get(LabId): Fetch (part 1)
                     
                     
                     
                     // Lab m5_get(LabId): Fetch (part 2)
                     
                     
               
                     // Lab m5_get(LabId): Instruction Types Decode and Immediate Decode
                     //_@1
                        // Types
                        assign FpgaPins_Fpga_CPU_is_i_instr_a1 = FpgaPins_Fpga_CPU_instr_a1[6:3] == 4'b0000 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b00100 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b00110 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b11001 ;
               
                        assign FpgaPins_Fpga_CPU_is_r_instr_a1 = FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b01011 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b01100 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b01110 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b10100 ;
               
                        assign FpgaPins_Fpga_CPU_is_s_instr_a1 = FpgaPins_Fpga_CPU_instr_a1[6:3] == 4'b0100;
               
                        assign FpgaPins_Fpga_CPU_is_b_instr_a1 = FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b11000;
               
                        assign FpgaPins_Fpga_CPU_is_j_instr_a1 = FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b11011;
               
                        assign FpgaPins_Fpga_CPU_is_u_instr_a1 = FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b00101 ||
                                      FpgaPins_Fpga_CPU_instr_a1[6:2] == 5'b01101;
                     
               
                     // Lab m5_get(LabId): Instruction Immediate Value Decoded
               
                        // Immediate
                        assign FpgaPins_Fpga_CPU_imm_a1[31:0]  =  FpgaPins_Fpga_CPU_is_i_instr_a1 ? {{21{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[30:20]} :
                                       FpgaPins_Fpga_CPU_is_s_instr_a1 ? {{21{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[30:25], FpgaPins_Fpga_CPU_instr_a1[11:7]} :
                                       FpgaPins_Fpga_CPU_is_b_instr_a1 ? {{20{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[7], FpgaPins_Fpga_CPU_instr_a1[30:25], FpgaPins_Fpga_CPU_instr_a1[11:8], 1'b0} :
                                       FpgaPins_Fpga_CPU_is_u_instr_a1 ? {FpgaPins_Fpga_CPU_instr_a1[31:12], 12'b0} :
                                       FpgaPins_Fpga_CPU_is_j_instr_a1 ? {{12{FpgaPins_Fpga_CPU_instr_a1[31]}}, FpgaPins_Fpga_CPU_instr_a1[19:12], FpgaPins_Fpga_CPU_instr_a1[20], FpgaPins_Fpga_CPU_instr_a1[30:21], 1'b0} :
                                                      32'b0 ;
                     
               
                     
                     // Lab m5_get(LabId): Instruction Immediate Valid
                     
                     
               
                     // Lab m5_get(LabId): Instruction Field Decode
                     
                     //_@1
                        assign FpgaPins_Fpga_CPU_funct7_valid_a1 = FpgaPins_Fpga_CPU_is_r_instr_a1;
                        assign FpgaPins_Fpga_CPU_funct3_valid_a1 = FpgaPins_Fpga_CPU_is_r_instr_a1 || FpgaPins_Fpga_CPU_is_i_instr_a1 || FpgaPins_Fpga_CPU_is_s_instr_a1 || FpgaPins_Fpga_CPU_is_b_instr_a1;
                        assign FpgaPins_Fpga_CPU_rs1_valid_a1    = FpgaPins_Fpga_CPU_is_r_instr_a1 || FpgaPins_Fpga_CPU_is_i_instr_a1 || FpgaPins_Fpga_CPU_is_s_instr_a1 || FpgaPins_Fpga_CPU_is_b_instr_a1;
                        assign FpgaPins_Fpga_CPU_rs2_valid_a1    = FpgaPins_Fpga_CPU_is_r_instr_a1 || FpgaPins_Fpga_CPU_is_s_instr_a1 || FpgaPins_Fpga_CPU_is_b_instr_a1 ;
                        assign FpgaPins_Fpga_CPU_rd_valid_a1     = FpgaPins_Fpga_CPU_is_r_instr_a1 || FpgaPins_Fpga_CPU_is_i_instr_a1 || FpgaPins_Fpga_CPU_is_u_instr_a1 || FpgaPins_Fpga_CPU_is_j_instr_a1;
                     
               
                     
                     // Lab m5_get(LabId): Instruction Decode
                     
                     
                     
               
                     
                     
                     
                     // Lab m5_get(LabId): Register File Read
                     
                     
                     
                     
                     
                     
               
                     
                     
                     // Lab m5_get(LabId): Register File Read (part 2)
                     
                     
               
                     
                     // Lab m5_get(LabId): Arithmetic Logic Unit
                     
                     
                     
               
                     // Lab m5_get(LabId): Register File Write
                     
                     
               
                     
                     // Lab m5_get(LabId): Branches (part 1)
                     
                     
                     
               
                     
                     // Lab m5_get(LabId): Branches (part 2)
                     
                     
                     
                     
               
                     
                     // Lab m5_get(LabId): Testbench
                     
                     
               
                     
                     // Lab m5_get(LabId): 3-Cycle Valid
                     
                     
               
                     // Lab m5_get(LabId): 3-Cycle RISC-V (part 1)
                     
                     
                     //_@1
                        assign FpgaPins_Fpga_CPU_inc_pc_a1[31:0] = FpgaPins_Fpga_CPU_pc_a1 + 32'd4;
                     //_@3
                        assign FpgaPins_Fpga_CPU_valid_taken_br_a3 = FpgaPins_Fpga_CPU_valid_a3 && FpgaPins_Fpga_CPU_taken_br_a3;
                     
               
                     // Lab m5_get(LabId): 3-Cycle RISC-V (part 2)
                     
                     
                     
                     
                     
                     
               
                     // Lab m5_get(LabId): Register File Bypass
                     
                     
               
                     // Lab m5_get(LabId): Determining Branch Shadow
                     
                     
                     
               
                     // Lab m5_get(LabId): Complete Instruction Decode
                     
                     //_@1
                        assign FpgaPins_Fpga_CPU_is_lui_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[6:0] ==        7'b0110111 ;
                        assign FpgaPins_Fpga_CPU_is_auipc_a1   =  FpgaPins_Fpga_CPU_dec_bits_a1[6:0] ==        7'b0010111 ;
                        assign FpgaPins_Fpga_CPU_is_jal_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[6:0] ==        7'b1101111 ;
                        assign FpgaPins_Fpga_CPU_is_jalr_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b000_1100111 ;
               
                        assign FpgaPins_Fpga_CPU_is_load_a1    =  FpgaPins_Fpga_CPU_opcode_a1        ==        7'b0000011 ;
               
                        //$is_sb      =  $dec_bits[9:0] ==   10'b000_0100011 ;
                        //$is_sh      =  $dec_bits[9:0] ==   10'b001_0100011 ;
                        //$is_sw      =  $dec_bits[9:0] ==   10'b010_0100011 ;
               
                        assign FpgaPins_Fpga_CPU_is_slti_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b010_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_sltiu_a1   =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b011_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_xori_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b100_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_ori_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b110_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_andi_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b111_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_slli_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_001_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_srli_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_101_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_srai_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b1_101_0010011 ;
               
                        assign FpgaPins_Fpga_CPU_is_sub_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b1_000_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_sll_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_001_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_slt_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_010_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_sltu_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_011_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_xor_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_100_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_srl_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_101_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_sra_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b1_101_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_or_a1      =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_110_0110011 ;
                        assign FpgaPins_Fpga_CPU_is_and_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_111_0110011 ;
               
                     
               
                     // Lab m5_get(LabId): Complete ALU
                     
                     //_@3
                        /* verilator lint_off WIDTH */
                        assign FpgaPins_Fpga_CPU_sltu_rslt_a3[31:0]      =   FpgaPins_Fpga_CPU_src1_value_a3 < FpgaPins_Fpga_CPU_src2_value_a3 ;
                        assign FpgaPins_Fpga_CPU_sltiu_rslt_a3[31:0]     =   FpgaPins_Fpga_CPU_src1_value_a3 < FpgaPins_Fpga_CPU_imm_a3;
                        /* verilator lint_on WIDTH */
                     
               
                     // Lab m5_get(LabId): Redirect Loads
                     
                     
                     //_@3
                        assign FpgaPins_Fpga_CPU_valid_load_a3 = FpgaPins_Fpga_CPU_valid_a3 && FpgaPins_Fpga_CPU_is_load_a3;
                     
               
                     // Lab m5_get(LabId): Load Data
                     
                     
                     
               
                     // Lab m5_get(LabId): Data Memory
                     //_@4
                        assign FpgaPins_Fpga_CPU_dmem_wr_en_a4          = FpgaPins_Fpga_CPU_is_s_instr_a4 && FpgaPins_Fpga_CPU_valid_a4;
                        assign FpgaPins_Fpga_CPU_dmem_wr_data_a4[31:0]  = FpgaPins_Fpga_CPU_src2_value_a4;
                        assign FpgaPins_Fpga_CPU_dmem_rd_en_a4          = FpgaPins_Fpga_CPU_is_load_a4;
                        assign FpgaPins_Fpga_CPU_dmem_addr_a4[2:0]      = FpgaPins_Fpga_CPU_result_a4[4:2];
               
                     //_@5
                        assign FpgaPins_Fpga_CPU_ld_data_a5[31:0]       = FpgaPins_Fpga_CPU_dmem_rd_data_a5;
               
                     //_\source /raw.githubusercontent.com/stevehoover/MESTCourse/main/tlvlib/riscvshelllib.tlv 50   // Instantiated from top.tlv, 504 as: m4+dmem(@4)
                        // Data Memory
                        //_@4
                           for (dmem = 0; dmem <= 7; dmem++) begin : L1_FpgaPins_Fpga_CPU_Dmem //_/dmem

                              // For $wr.
                              logic L1_wr_a4;

                              assign L1_wr_a4 = FpgaPins_Fpga_CPU_dmem_wr_en_a4 && (FpgaPins_Fpga_CPU_dmem_addr_a4[2:0] == dmem);
                              assign FpgaPins_Fpga_CPU_Dmem_value_a4[dmem][31:0] = FpgaPins_Fpga_CPU_reset_a4 ?   dmem :
                                             L1_wr_a4        ?   FpgaPins_Fpga_CPU_dmem_wr_data_a4 :
                                                            FpgaPins_Fpga_CPU_Dmem_value_a5[dmem][31:0];
                           end
                     
                           //_?$dmem_rd_en
                              assign FpgaPins_Fpga_CPU_dmem_rd_data_a4[31:0] = FpgaPins_Fpga_CPU_Dmem_value_a5[FpgaPins_Fpga_CPU_dmem_addr_a4[2:0]];
                           `BOGUS_USE(FpgaPins_Fpga_CPU_dmem_rd_data_a4)
                     //_\end_source
                     
               
                  // Lab m5_get(LabId): Load/Store in Program
               
                  //_|cpu
                     
                  
               
                     // Lab m5_get(LabId): Jumps
                     
                     
               
                     //_@3
                        assign FpgaPins_Fpga_CPU_is_jump_a3    =  FpgaPins_Fpga_CPU_is_jal_a3 || FpgaPins_Fpga_CPU_is_jalr_a3;
                        assign FpgaPins_Fpga_CPU_jalr_tgt_pc_a3[31:0]   =  FpgaPins_Fpga_CPU_src1_value_a3 + FpgaPins_Fpga_CPU_imm_a3;
                        assign FpgaPins_Fpga_CPU_valid_jump_a3 =  FpgaPins_Fpga_CPU_is_jump_a3 && FpgaPins_Fpga_CPU_valid_a3;
                     
               
               
               
                     // Logic that changes throughout.
               
               
                     //_@0
                     
                        
                                                      
                     
                        
                                       
                                                         
                     
                        
                                       
                                                               
                     
                        
                                       
                                                               
                     
                        
                                       
                                       
                                                               
                     
                        assign FpgaPins_Fpga_CPU_pc_a0[31:0]   =  FpgaPins_Fpga_CPU_reset_a1                     ?  '0 :
                                       FpgaPins_Fpga_CPU_valid_taken_br_a3            ?  FpgaPins_Fpga_CPU_br_tgt_pc_a3   :
                                       FpgaPins_Fpga_CPU_valid_load_a3                ?  FpgaPins_Fpga_CPU_inc_pc_a3      :
                                       FpgaPins_Fpga_CPU_valid_jump_a3 && FpgaPins_Fpga_CPU_is_jal_a3  ?  FpgaPins_Fpga_CPU_br_tgt_pc_a3   :
                                       FpgaPins_Fpga_CPU_valid_jump_a3 && FpgaPins_Fpga_CPU_is_jalr_a3 ?  FpgaPins_Fpga_CPU_jalr_tgt_pc_a3 :
                                                                        FpgaPins_Fpga_CPU_inc_pc_a1 ;
                     
               
                     
                     //_@2
                        assign FpgaPins_Fpga_CPU_br_tgt_pc_a2[31:0] = FpgaPins_Fpga_CPU_pc_a2 + FpgaPins_Fpga_CPU_imm_a2;
                     
               
                     
                     //_@0
                        assign FpgaPins_Fpga_CPU_imem_rd_en_a0                          = !FpgaPins_Fpga_CPU_reset_a0;
                        assign FpgaPins_Fpga_CPU_imem_rd_addr_a0[4-1:0] = FpgaPins_Fpga_CPU_pc_a0[4+1:2];
                     //_@1
                        assign FpgaPins_Fpga_CPU_instr_a1[31:0]                         = FpgaPins_Fpga_CPU_imem_rd_data_a1[31:0];
                        //`BOGUS_USE($instr)
                     
               
                     
                     
                        
                        
                        
                        
                        
                        
                        
                              // Other fields
                     //_@1
                        //_?$funct7_valid
                           assign FpgaPins_Fpga_CPU_funct7_a1[6:0] = FpgaPins_Fpga_CPU_instr_a1[31:25];
                        //_?$funct3_valid
                           assign FpgaPins_Fpga_CPU_funct3_a1[2:0] = FpgaPins_Fpga_CPU_instr_a1[14:12];
                        //_?$rs1_valid
                           assign FpgaPins_Fpga_CPU_rs1_a1[4:0]    = FpgaPins_Fpga_CPU_instr_a1[19:15];
                        //_?$rs2_valid
                           assign FpgaPins_Fpga_CPU_rs2_a1[4:0]    = FpgaPins_Fpga_CPU_instr_a1[24:20];
                        //_?$rd_valid
                           assign FpgaPins_Fpga_CPU_rd_a1[4:0]     = FpgaPins_Fpga_CPU_instr_a1[11:7];
                        assign FpgaPins_Fpga_CPU_opcode_a1[6:0]    = FpgaPins_Fpga_CPU_instr_a1[6:0];
                        //`BOGUS_USE($funct7 $funct3 $opcode $funct3)
                     
               
                     
                     //_@1
                        assign FpgaPins_Fpga_CPU_dec_bits_a1[10:0] = {FpgaPins_Fpga_CPU_funct7_a1[5], FpgaPins_Fpga_CPU_funct3_a1, FpgaPins_Fpga_CPU_opcode_a1};
                        assign FpgaPins_Fpga_CPU_is_beq_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b000_1100011 ;
                        assign FpgaPins_Fpga_CPU_is_bne_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b001_1100011 ;
                        assign FpgaPins_Fpga_CPU_is_blt_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b100_1100011 ;
                        assign FpgaPins_Fpga_CPU_is_bge_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b101_1100011 ;
                        assign FpgaPins_Fpga_CPU_is_bltu_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b110_1100011 ;
                        assign FpgaPins_Fpga_CPU_is_bgeu_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b111_1100011 ;
               
                        assign FpgaPins_Fpga_CPU_is_addi_a1    =  FpgaPins_Fpga_CPU_dec_bits_a1[9:0] ==   10'b000_0010011 ;
                        assign FpgaPins_Fpga_CPU_is_add_a1     =  FpgaPins_Fpga_CPU_dec_bits_a1      == 11'b0_000_0110011 ;
                     
               
                     //_@2
                     
                        assign FpgaPins_Fpga_CPU_rf_rd_en1_a2           =  FpgaPins_Fpga_CPU_rs1_valid_a2;
                        assign FpgaPins_Fpga_CPU_rf_rd_en2_a2           =  FpgaPins_Fpga_CPU_rs2_valid_a2;
                        assign FpgaPins_Fpga_CPU_rf_rd_index1_a2[4:0]   =  FpgaPins_Fpga_CPU_rs1_a2;
                        assign FpgaPins_Fpga_CPU_rf_rd_index2_a2[4:0]   =  FpgaPins_Fpga_CPU_rs2_a2;
                     
               
                     
                     
                     
                        
                        
                     
                     
                        assign FpgaPins_Fpga_CPU_src1_value_a2[31:0] =
                             (FpgaPins_Fpga_CPU_rf_wr_index_a3 == FpgaPins_Fpga_CPU_rf_rd_index1_a2) && FpgaPins_Fpga_CPU_rf_wr_en_a3
                                 ?  FpgaPins_Fpga_CPU_result_a3   :
                                    FpgaPins_Fpga_CPU_rf_rd_data1_a2 ;
                        assign FpgaPins_Fpga_CPU_src2_value_a2[31:0] =
                             (FpgaPins_Fpga_CPU_rf_wr_index_a3 == FpgaPins_Fpga_CPU_rf_rd_index2_a2) && FpgaPins_Fpga_CPU_rf_wr_en_a3
                                 ?  FpgaPins_Fpga_CPU_result_a3   :
                                    FpgaPins_Fpga_CPU_rf_rd_data2_a2 ;
                     
                     
               
                     //_@3
                     
                        
                        
                        
                     
                        
                        
                        
                     
                        
                        
                        
                     
                        assign FpgaPins_Fpga_CPU_rf_wr_en_a3            =  (FpgaPins_Fpga_CPU_rd_valid_a3 && FpgaPins_Fpga_CPU_valid_a3 && FpgaPins_Fpga_CPU_rd_a3 != 5'b0) || FpgaPins_Fpga_CPU_valid_load_a5;
                        assign FpgaPins_Fpga_CPU_rf_wr_index_a3[4:0]    =  FpgaPins_Fpga_CPU_valid_load_a5 ? FpgaPins_Fpga_CPU_rd_a5 : FpgaPins_Fpga_CPU_rd_a3;
                        assign FpgaPins_Fpga_CPU_rf_wr_data_a3[31:0]    =  FpgaPins_Fpga_CPU_valid_load_a5 ? FpgaPins_Fpga_CPU_ld_data_a5 : FpgaPins_Fpga_CPU_result_a3;
                     
               
                     /* verilator lint_off WIDTH */
               
                     
                     
                        
                                          
                                                      
                     
                     //_@3
                        assign FpgaPins_Fpga_CPU_result_a3[31:0] =   FpgaPins_Fpga_CPU_is_andi_a3    ?  FpgaPins_Fpga_CPU_src1_value_a3 & FpgaPins_Fpga_CPU_imm_a3 :
                                          FpgaPins_Fpga_CPU_is_ori_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 | FpgaPins_Fpga_CPU_imm_a3 :
                                          FpgaPins_Fpga_CPU_is_xori_a3    ?  FpgaPins_Fpga_CPU_src1_value_a3 ^ FpgaPins_Fpga_CPU_imm_a3 :
                                          (FpgaPins_Fpga_CPU_is_addi_a3 || FpgaPins_Fpga_CPU_is_load_a3 || FpgaPins_Fpga_CPU_is_s_instr_a3) ?  FpgaPins_Fpga_CPU_src1_value_a3 + FpgaPins_Fpga_CPU_imm_a3 :
                                          FpgaPins_Fpga_CPU_is_slli_a3    ?  FpgaPins_Fpga_CPU_src1_value_a3 << FpgaPins_Fpga_CPU_imm_a3[5:0]  :
                                          FpgaPins_Fpga_CPU_is_srli_a3    ?  FpgaPins_Fpga_CPU_src1_value_a3 >> FpgaPins_Fpga_CPU_imm_a3[5:0]  :
                                          FpgaPins_Fpga_CPU_is_and_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 & FpgaPins_Fpga_CPU_src2_value_a3 :
                                          FpgaPins_Fpga_CPU_is_or_a3      ?  FpgaPins_Fpga_CPU_src1_value_a3 | FpgaPins_Fpga_CPU_src2_value_a3 :
                                          FpgaPins_Fpga_CPU_is_xor_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 ^ FpgaPins_Fpga_CPU_src2_value_a3 :
                                          FpgaPins_Fpga_CPU_is_add_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 + FpgaPins_Fpga_CPU_src2_value_a3 :
                                          FpgaPins_Fpga_CPU_is_sub_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 - FpgaPins_Fpga_CPU_src2_value_a3 :
                                          FpgaPins_Fpga_CPU_is_sll_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 << FpgaPins_Fpga_CPU_src2_value_a3[4:0] :
                                          FpgaPins_Fpga_CPU_is_srl_a3     ?  FpgaPins_Fpga_CPU_src1_value_a3 >> FpgaPins_Fpga_CPU_src2_value_a3[4:0] :
                                          FpgaPins_Fpga_CPU_is_sltu_a3    ?  FpgaPins_Fpga_CPU_sltu_rslt_a3 :
                                          FpgaPins_Fpga_CPU_is_sltiu_a3   ?  FpgaPins_Fpga_CPU_sltiu_rslt_a3 :
                                          FpgaPins_Fpga_CPU_is_lui_a3     ?  {FpgaPins_Fpga_CPU_imm_a3[31:12], 12'b0} :
                                          FpgaPins_Fpga_CPU_is_auipc_a3   ?  FpgaPins_Fpga_CPU_pc_a3 + FpgaPins_Fpga_CPU_imm_a3 :
                                          FpgaPins_Fpga_CPU_is_jal_a3     ?  FpgaPins_Fpga_CPU_pc_a3 + 32'd4 :
                                          FpgaPins_Fpga_CPU_is_jalr_a3    ?  FpgaPins_Fpga_CPU_pc_a3 + 32'd4 :
                                          FpgaPins_Fpga_CPU_is_srai_a3    ?  {{32{FpgaPins_Fpga_CPU_src1_value_a3[31]}}, FpgaPins_Fpga_CPU_src1_value_a3} >> FpgaPins_Fpga_CPU_imm_a3[4:0] :
                                          FpgaPins_Fpga_CPU_is_slt_a3     ?  ((FpgaPins_Fpga_CPU_src1_value_a3[31] == FpgaPins_Fpga_CPU_src2_value_a3[31]) ? FpgaPins_Fpga_CPU_sltu_rslt_a3  : {31'b0, FpgaPins_Fpga_CPU_src1_value_a3[31]}) :
                                          FpgaPins_Fpga_CPU_is_slti_a3    ?  ((FpgaPins_Fpga_CPU_src1_value_a3[31] == FpgaPins_Fpga_CPU_imm_a3[31])        ? FpgaPins_Fpga_CPU_sltiu_rslt_a3 : {31'b0, FpgaPins_Fpga_CPU_src1_value_a3[31]}) :
                                          FpgaPins_Fpga_CPU_is_sra_a3     ?  {{32{FpgaPins_Fpga_CPU_src1_value_a3[31]}}, FpgaPins_Fpga_CPU_src1_value_a3} >> FpgaPins_Fpga_CPU_src2_value_a3[4:0] :
                                                         32'bx;
                     
               
                     /* verilator lint_on WIDTH */
               
                     
                     //_@3
                        assign FpgaPins_Fpga_CPU_taken_br_a3   =  FpgaPins_Fpga_CPU_is_beq_a3  ? (FpgaPins_Fpga_CPU_src1_value_a3 == FpgaPins_Fpga_CPU_src2_value_a3) :
                                       FpgaPins_Fpga_CPU_is_bne_a3  ? (FpgaPins_Fpga_CPU_src1_value_a3 != FpgaPins_Fpga_CPU_src2_value_a3) :
                                       FpgaPins_Fpga_CPU_is_blt_a3  ? ((FpgaPins_Fpga_CPU_src1_value_a3 < FpgaPins_Fpga_CPU_src2_value_a3)  ^ (FpgaPins_Fpga_CPU_src1_value_a3[31] != FpgaPins_Fpga_CPU_src2_value_a3[31])) :
                                       FpgaPins_Fpga_CPU_is_bge_a3  ? ((FpgaPins_Fpga_CPU_src1_value_a3 >= FpgaPins_Fpga_CPU_src2_value_a3) ^ (FpgaPins_Fpga_CPU_src1_value_a3[31] != FpgaPins_Fpga_CPU_src2_value_a3[31])) :
                                       FpgaPins_Fpga_CPU_is_bltu_a3 ? (FpgaPins_Fpga_CPU_src1_value_a3 < FpgaPins_Fpga_CPU_src2_value_a3)  :
                                       FpgaPins_Fpga_CPU_is_bgeu_a3 ? (FpgaPins_Fpga_CPU_src1_value_a3 >= FpgaPins_Fpga_CPU_src2_value_a3) :
                                                  1'b0;
                        //`BOGUS_USE($taken_br)
                     
               
                     
                     
                        
                        
                                 
                                          
                     
                     
                        
                     
                     
                        
                                   
                     
                     //_@3
                        assign FpgaPins_Fpga_CPU_valid_a3 = !(FpgaPins_Fpga_CPU_valid_taken_br_a4 || FpgaPins_Fpga_CPU_valid_taken_br_a5 ||
                                   FpgaPins_Fpga_CPU_valid_load_a4     || FpgaPins_Fpga_CPU_valid_load_a5     ||
                                   FpgaPins_Fpga_CPU_valid_jump_a4     || FpgaPins_Fpga_CPU_valid_jump_a5);
                     
               
                     //_@1
                        
                        
                        
                        assign passed = FpgaPins_Fpga_CPU_Xreg_value_a6[15] == (1+2+3+4+5+6+7+8+9);
                        
                        
                        
               
               
                  assign failed = 1'b0;
               
                  //_|cpu
                     
                     // IMem
                     //_\source /raw.githubusercontent.com/stevehoover/MESTCourse/main/tlvlib/riscvshelllib.tlv 18   // Instantiated from top.tlv, 740 as: m4+imem(@1)
                        // Instruction Memory containing program.
                        //_@1
                           /*SV_plus*/
                              // The program in an instruction memory.
                              logic [31:0] instrs [0:10-1];
                              assign instrs[0] = {7'b0000000, 5'd0, 5'd0, 3'b000, 5'd10, 7'b0110011}; assign instrs[1] = {7'b0000000, 5'd0, 5'd10, 3'b000, 5'd14, 7'b0110011}; assign instrs[2] = {12'b000000001010, 5'd10, 3'b000, 5'd12, 7'b0010011}; assign instrs[3] = {7'b0000000, 5'd0, 5'd10, 3'b000, 5'd13, 7'b0110011}; assign instrs[4] = {7'b0000000, 5'd14, 5'd13, 3'b000, 5'd14, 7'b0110011}; assign instrs[5] = {12'b000000000001, 5'd13, 3'b000, 5'd13, 7'b0010011}; assign instrs[6] = {1'b1, 6'b111111, 5'd12, 5'd13, 3'b100, 4'b1100, 1'b1, 7'b1100011}; assign instrs[7] = {7'b0000000, 5'd0, 5'd14, 3'b000, 5'd10, 7'b0110011}; assign instrs[8] = {7'b0000000, 5'd10, 5'd0, 3'b010, 5'b00100, 7'b0100011}; assign instrs[9] = {12'b000000000100, 5'd0, 3'b010, 5'd15, 7'b0000011}; 
                           for (imem = 0; imem <= 9; imem++) begin : L1_FpgaPins_Fpga_CPU_Imem //_/imem
                              assign FpgaPins_Fpga_CPU_Imem_instr_a1[imem][31:0] = instrs[imem];
                           end
                           //_?$imem_rd_en
                              assign FpgaPins_Fpga_CPU_imem_rd_data_a1[31:0] = FpgaPins_Fpga_CPU_Imem_instr_a1[FpgaPins_Fpga_CPU_imem_rd_addr_a1];
                     //_\end_source    // Args: (read stage)
                     
               
                     // Args: (read stage, write stage) - if equal, no register bypass is required
                     
                     //_\source /raw.githubusercontent.com/stevehoover/MESTCourse/main/tlvlib/riscvshelllib.tlv 33   // Instantiated from top.tlv, 745 as: m4+rf(m5_get(rf_rd_stage), m5_get(rf_wr_stage))
                        // Reg File
                        //_@3
                           for (xreg = 0; xreg <= 15; xreg++) begin : L1_FpgaPins_Fpga_CPU_Xreg //_/xreg

                              // For $wr.
                              logic L1_wr_a3;

                              assign L1_wr_a3 = FpgaPins_Fpga_CPU_rf_wr_en_a3 && (FpgaPins_Fpga_CPU_rf_wr_index_a3 != 5'b0) && (FpgaPins_Fpga_CPU_rf_wr_index_a3 == xreg);
                              assign FpgaPins_Fpga_CPU_Xreg_value_a3[xreg][31:0] = FpgaPins_Fpga_CPU_reset_a3 ?   xreg           :
                                             L1_wr_a3        ?   FpgaPins_Fpga_CPU_rf_wr_data_a3 :
                                                            FpgaPins_Fpga_CPU_Xreg_value_a4[xreg][31:0];
                           end
                        //_@2
                           //_?$rf_rd_en1
                              assign FpgaPins_Fpga_CPU_rf_rd_data1_a2[31:0] = FpgaPins_Fpga_CPU_Xreg_value_a4[FpgaPins_Fpga_CPU_rf_rd_index1_a2[3:0]];
                           //_?$rf_rd_en2
                              assign FpgaPins_Fpga_CPU_rf_rd_data2_a2[31:0] = FpgaPins_Fpga_CPU_Xreg_value_a4[FpgaPins_Fpga_CPU_rf_rd_index2_a2[3:0]];
                           `BOGUS_USE(FpgaPins_Fpga_CPU_rf_rd_data1_a2 FpgaPins_Fpga_CPU_rf_rd_data2_a2)
                     //_\end_source
                     
               
                  // ============================================================================================================
               
                  // Connect Tiny Tapeout outputs.
                  // Note that my_design will be under /fpga_pins/fpga.
                  assign uo_out = {6'b0, failed, passed};
                  
                  
               
                      // For visualisation, argument should be at least equal to the last stage of CPU logic. @4 would work for all labs.
               //_\end_source
            
            //_\end_source
   
      // LEDs.
      
   
      // 7-Segment
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 395   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 346 as: m4+fpga_sseg.
         for (digit = 0; digit <= 0; digit++) begin : L1_Digit //_/digit
            
            for (leds = 0; leds <= 7; leds++) begin : L2_Leds //_/leds

               // For $viz_lit.
               logic L2_viz_lit_a0;

               assign L2_viz_lit_a0 = (! L0_sseg_digit_n_a0[digit]) && ! ((leds == 7) ? L0_sseg_decimal_point_n_a0 : L0_sseg_segment_n_a0[leds % 7]);
               
            end
         end
      //_\end_source
   
      // slideswitches
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 454   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 349 as: m4+fpga_switch.
         for (switch = 0; switch <= 7; switch++) begin : L1_Switch //_/switch

            // For $viz_switch.
            logic L1_viz_switch_a0;

            assign L1_viz_switch_a0 = L0_slideswitch_a0[switch];
            
         end
      //_\end_source
   
      // pushbuttons
      
   //_\end_source
   // Label the switch inputs [0..7] (1..8 on the physical switch panel) (top-to-bottom).
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/af18805ea79802b83477cf86aff503e97ed7394a/tlvlib/tinytapeoutlib.tlv 73   // Instantiated from top.tlv, 863 as: m5+tt_input_labels_viz(m5_get(input_labels))
      for (input_label = 0; input_label <= 7; input_label++) begin : L1_InputLabel //_/input_label
         
      end
   //_\end_source

//_\SV
endmodule


// Undefine macros defined by SandPiper.
`undef BOGUS_USE
